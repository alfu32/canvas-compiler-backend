module utils



pub struct Ref {
	pub mut:
	ref string
}
