module entities
