module entities

